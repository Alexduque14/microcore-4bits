module bcd_display(
	input wire [3:0] in,
	output reg [6:0] disp
);

always @(*) begin
	case (in) 			
		4'b0000: disp = 7'b0000001;	//0
		4'b0001: disp = 7'b1001111;	//1
		4'b0010: disp = 7'b0010010;	//2
		4'b0011: disp = 7'b0000110;	//3
		4'b0100: disp = 7'b1001100;	//4
		4'b0101: disp = 7'b0100100;	//5
		4'b0110: disp = 7'b0100000;	//6
		4'b0111:	disp = 7'b0001111;	//7
		4'b1000:	disp = 7'b0000000;	//8
		4'b1001:	disp = 7'b0000100;	//9
		4'b1010:	disp = 7'b0001000; 	//10(A)
		4'b1011:	disp = 7'b1100000;	//11(b)
		4'b1100:	disp = 7'b0110001;	//12(C)
		4'b1101:	disp = 7'b1000010;	//13(d)
		4'b1110:	disp = 7'b0110000;	//14(E)
		4'b1111:	disp = 7'b0111000;	//15(F)
		default: disp = 7'b1111111;	//off
		endcase
	end
endmodule
		